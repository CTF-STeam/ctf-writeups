module check(
    input clk,

    input [6:0] data,
    output wire open_safe
);

reg [6:0] memory [7:0];
reg [2:0] idx = 0;

wire [55:0] magic = {
    {memory[0], memory[5]},
    {memory[6], memory[2]},
    {memory[4], memory[3]},
    {memory[7], memory[1]}
};

wire [55:0] kittens = { magic[9:0],  magic[41:22], magic[21:10], magic[55:42] };
assign open_safe = kittens == 56'd3008192072309708;

always_ff @(posedge clk) begin
    memory[idx] <= data;
    idx <= idx + 5;
end

endmodule

/*
kittens
00001010101011111110111101001011111000101101101111001100
0000101010 10111111101111010010 111110001011 01101111001100
9        0 41                22 21        10 55          42

magic
01101111001100 10111111101111010010 111110001011 0000101010
55          42 41                22 21        10 9        0
01101111001100101111111011110100101111100010110000101010

0110111 1001100 1011111 1101111 0100101 1111000 1011000 0101010
      0       5       6       2       4       3       7       1

memory

1011000 1011111 1001100 0100101 1111000 1101111 0101010 0110111
      7       6       5       4       3       2       1       0

0000101 1001100 1101111 1010010 1110111 0101111 1000101 0110111
      0       1       2       3       4       5       6       7

data
0110111 1001100 1101111 1011000 0100101 0101010 1011111 1111000
      0       5       2       7       4       1       6       3

00110111 01001100 01101111 01011000 00100101 00101010 01011111 01111000
7LoX%*_x

*/

